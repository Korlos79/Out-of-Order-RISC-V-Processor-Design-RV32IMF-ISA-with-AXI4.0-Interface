module alu (
    input  wire        clk,
    input  wire        rst_n,
    input  wire [31:0] A,
    input  wire [31:0] B,
    input  wire [6:0]  opcode,
    input  wire [2:0]  branch,
    
    // --- OUTPUTS ĐƯỢC TÁCH BIỆT ---
    output reg  [31:0] alu_result,    // Kết quả cơ bản (ADD, SUB...) - Có ngay
    output wire [31:0] md_result,     // Kết quả Nhân/Chia - Có trễ
    output wire        md_busy,       // Trạng thái bận của khối Nhân/Chia
    output wire        md_done,       // Báo xong của khối Nhân/Chia
    
    output reg         Z
);

    // --- 1. DEFINITIONS ---
    localparam beq  = 3'b000;
    localparam bne  = 3'b001;
    localparam blt  = 3'b100;
    localparam bge  = 3'b101;
    localparam bltu = 3'b110;
    localparam bgeu = 3'b111;

    // --- 2. M-EXTENSION HANDLING ---
    wire is_m_op = (opcode >= 6'd9 && opcode <= 6'd16);

    reg [4:0] muldiv_op_sel;
    always @(*) begin
        if (is_m_op) 
            muldiv_op_sel = 6'b010000 + (opcode - 6'd9);
        else 
            muldiv_op_sel = 6'b00000;
    end

    // Instantiate M-Extension Unit
    // Kết quả nối thẳng ra output md_result, md_busy, md_done
    rv32m_muldiv_split U_MULDIV (
        .clk(clk),
        .rst_n(rst_n),
        .op_valid(is_m_op),     
        .op_sel(muldiv_op_sel),
        .rs1(A),
        .rs2(B),
        .busy(md_busy),
        .done(md_done),
        .result(md_result)
    );

    // --- 3. BASE INTEGER ALU LOGIC ---
    // Logic tổ hợp, luôn tính toán dựa trên A, B và Opcode hiện tại
    always @(*) begin
        case(opcode)
            6'd0: alu_result = A + B;             // ADD
            6'd1: alu_result = A << B[4:0];       // SLL
            6'd2: alu_result = ($signed(A) < $signed(B)) ? 32'd1 : 32'd0;     // SLT
            6'd3: alu_result = ($unsigned(A) < $unsigned(B)) ? 32'd1 : 32'd0; // SLTU
            6'd4: alu_result = A ^ B;             // XOR
            6'd5: alu_result = A >> B[4:0];       // SRL
            6'd6: alu_result = A | B;             // OR
            6'd7: alu_result = A & B;             // AND
            6'd8: alu_result = A - B;             // SUB
            6'd17: alu_result = $signed(A) >>> B[4:0]; // SRA (Thêm lệnh này)
            default: alu_result = 32'd0;
        endcase
    end

    // --- 4. BRANCH COMPARATOR ---
    always @(*) begin
        case (branch)
            beq:  Z = (A == B);
            bne:  Z = (A != B);
            blt:  Z = ($signed(A) < $signed(B));
            bge:  Z = ($signed(A) >= $signed(B)); 
            bltu: Z = ($unsigned(A) < $unsigned(B));
            bgeu: Z = ($unsigned(A) >= $unsigned(B));
            default: Z = 1'b0;
        endcase
    end

endmodule