`timescale 1ns / 1ps

module tb_iter_mul32();

    // --- 1. Signal Declaration ---
    reg clk;
    reg rst_n;
    reg start;
    reg [4:0] op_sel;
    reg [31:0] rs1;
    reg [31:0] rs2;

    wire busy;
    wire done;
    wire [31:0] result;

    // --- 2. Opcodes (Local Copy for TB) ---
    localparam OP_MUL    = 5'b10000;
    localparam OP_MULH   = 5'b10001; // Signed x Signed (High)
    localparam OP_MULHSU = 5'b10010; // Signed x Unsigned (High)
    localparam OP_MULHU  = 5'b10011; // Unsigned x Unsigned (High)

    // --- 3. Instantiate DUT ---
    iter_mul32 uut (
        .clk(clk),
        .rst_n(rst_n),
        .start(start),
        .op_sel(op_sel),
        .rs1(rs1),
        .rs2(rs2),
        .busy(busy),
        .done(done),
        .result(result)
    );

    // --- 4. Clock Generation (100MHz) ---
    always #5 clk = ~clk;

    // --- 5. Monitor Output ---
    // Hiển thị kết quả ngay khi 'done' bật lên (trễ 4 chu kì so với input)
    integer output_cnt = 0;
	 real    start_time;
    always @(posedge clk) begin
        if (done) begin
            output_cnt = output_cnt + 1;
            $display("[OUTPUT %0d] Time %t | Cycle %0d | Result = %h (%0d)", output_cnt, $time, ($realtime - start_time)/10 - 1, result, $signed(result));
        end
    end

    // --- 6. Task: Gửi lệnh (Send Command) ---
    task send_cmd;
        input [4:0] opcode;
        input [31:0] in1;
        input [31:0] in2;
        input [127:0] comment; // Chuỗi ký tự mô tả
        begin
            @(posedge clk); // Đợi cạnh lên để đồng bộ
            start  <= 1;
				start_time = $realtime;
            op_sel <= opcode;
            rs1    <= in1;
            rs2    <= in2;
            
            $display("[INPUT]  Time %t | %s | RS1=%h (%0d), RS2=%h (%0d)", 
                     $time, comment, in1, $signed(in1), in2, $signed(in2));
            
            @(posedge clk);
            start  <= 0; // Tắt start sau 1 chu kì (tạo xung pulse)
            // Lưu ý: Task này tốn 1 chu kì clock để gửi xong 1 lệnh
        end
    endtask

    // --- 7. Main Test Sequence ---
    initial begin
        // Init
        clk = 0; rst_n = 0; start = 0;
        op_sel = 0; rs1 = 0; rs2 = 0;

        // Reset
        $display("=== RESET SYSTEM ===");
        #20 rst_n = 1;
        #20;

        // ============================================================
        // TEST CASE 1: Lệnh MUL (Lấy 32-bit thấp)
        // ============================================================
        $display("\n=== TEST 1: MUL (Low 32-bit) ===");
        
        // 10 * -5 = -50 (FFFF_FFCE)
        send_cmd(OP_MUL, 32'd10, -32'd5, "10 * -5");
        
        #50; // Đợi kết quả trôi ra hết

        // ============================================================
        // TEST CASE 2: Các lệnh High (MULH, MULHSU, MULHU)
        // ============================================================
        $display("\n=== TEST 2: High Part Multiplication ===");
        
        // Setup: A = -2 (FFFFFFFE), B = -2 (FFFFFFFE)
        // Tích 64-bit: (-2) * (-2) = 4 (00000000_00000004)
        
        // 2.1 MULH (Signed * Signed) -> High part = 0
        send_cmd(OP_MULH, -32'd2, -32'd2, "MULH (-2 * -2)");
        #50;

        // Setup: A = Max Int (7FFFFFFF), B = 2
        // Tích: 2 * (2^31 - 1) = 2^32 - 2 = 00000000_FFFFFFFE (High=0, Low=-2)
        // Nhưng nếu là MULH thì ta cần số lớn hơn để High != 0
        // Thử: MaxInt * MaxInt = ~ 2^62 (High sẽ rất lớn)
        send_cmd(OP_MULH, 32'h7FFFFFFF, 32'h7FFFFFFF, "MULH (Max * Max)");
        #50;

        // ============================================================
        // TEST CASE 3: PIPELINE STRESS TEST (Back-to-back Inputs)
        // Gửi 3 lệnh liên tiếp không nghỉ
        // ============================================================
        $display("\n=== TEST 3: Pipeline Throughput (3 ops back-to-back) ===");
        
        // Chú ý: Vì task send_cmd đã có @(posedge clk) ở cuối để tắt start,
        // nên gọi liên tiếp các task này sẽ tạo ra chuỗi lệnh liên tục.
        
        // Op 1: 3 * 4 = 12
        send_cmd(OP_MUL, 32'd3, 32'd4, "Burst 1: 3 * 4");
        
        // Op 2: 5 * 6 = 30
        send_cmd(OP_MUL, 32'd5, 32'd6, "Burst 2: 5 * 6");
        
        // Op 3: 10 * 10 = 100
        send_cmd(OP_MUL, 32'd10, 32'd10, "Burst 3: 10 * 10");

        // Đợi kết quả
        #100;
        
        $display("\n=== END OF SIMULATION ===");
        $finish;
    end

endmodule