`timescale 1ns / 1ps

module tb_memory_system_full;

    // --- 1. Tín hiệu Clock & Reset ---
    reg clk;
    reg rst_n;

    // --- 2. Tín hiệu giả lập CPU -> IFU ---
    reg  [31:0] pc;
    wire [31:0] instr;
    wire        ifu_stall;

    // --- 3. Tín hiệu giả lập CPU -> LSU ---
    reg         lsu_we;     // Write Enable
    reg         lsu_re;     // Read Enable
    reg  [2:0]  lsu_mode;   // funct3
    reg  [31:0] lsu_addr;
    reg  [31:0] lsu_wdata;
    wire [31:0] lsu_rdata;
    wire        lsu_stall;

    // --- 4. Các dây nối AXI (Interconnect <-> Modules) ---
    // IFU -> Interconnect
    wire [31:0] ifu_araddr; wire ifu_arvalid, ifu_arready;
    wire [31:0] ifu_rdata;  wire ifu_rvalid, ifu_rready;

    // LSU -> Interconnect
    wire [31:0] lsu_awaddr; wire lsu_awvalid, lsu_awready;
    wire [31:0] lsu_wdata_wire; wire [3:0] lsu_wstrb; wire lsu_wvalid, lsu_wready;
    wire lsu_bvalid, lsu_bready;
    wire [31:0] lsu_araddr; wire lsu_arvalid, lsu_arready;
    wire [31:0] lsu_rdata_wire; wire lsu_rvalid, lsu_rready;

    // Interconnect -> RAM (Master Port)
    wire [31:0] mem_awaddr; wire mem_awvalid, mem_awready;
    wire [31:0] mem_wdata;  wire [3:0] mem_wstrb; wire mem_wvalid, mem_wready;
    wire mem_bvalid, mem_bready;
    wire [31:0] mem_araddr; wire mem_arvalid, mem_arready;
    wire [31:0] mem_rdata;  wire mem_rvalid, mem_rready;

    // =========================================================
    // INSTANTIATE CÁC MODULE (DUT)
    // =========================================================

    // 1. IFU (Instruction Fetch)
    instruction_Mem DUT_IFU (
        .clk(clk), .rst_n(rst_n),
        .addr(pc), .inst(instr), .stall_out(ifu_stall),
        // AXI Read Only
        .m_axi_araddr(ifu_araddr), .m_axi_arvalid(ifu_arvalid), .m_axi_arready(ifu_arready),
        .m_axi_rdata(ifu_rdata),   .m_axi_rvalid(ifu_rvalid),   .m_axi_rready(ifu_rready)
    );

    // 2. LSU (Load Store)
    dmem DUT_LSU (
        .clk(clk), .rst_n(rst_n),
        .we(lsu_we), .re(lsu_re), .mode(lsu_mode),
        .addr(lsu_addr), .write_data(lsu_wdata), .mem_out(lsu_rdata), .stall_out(lsu_stall),
        // AXI Write
        .m_axi_awaddr(lsu_awaddr), .m_axi_awvalid(lsu_awvalid), .m_axi_awready(lsu_awready),
        .m_axi_wdata(lsu_wdata_wire), .m_axi_wstrb(lsu_wstrb), .m_axi_wvalid(lsu_wvalid), .m_axi_wready(lsu_wready),
        .m_axi_bvalid(lsu_bvalid), .m_axi_bready(lsu_bready),
        // AXI Read
        .m_axi_araddr(lsu_araddr), .m_axi_arvalid(lsu_arvalid), .m_axi_arready(lsu_arready),
        .m_axi_rdata(lsu_rdata_wire), .m_axi_rvalid(lsu_rvalid), .m_axi_rready(lsu_rready)
    );

    // 3. INTERCONNECT (Trọng tài)
    axi4_interconnect_2x1 DUT_INTERCONNECT (
        .clk(clk), .rst_n(rst_n),
        
        // Slave 0: IFU
        .s0_axi_araddr(ifu_araddr), .s0_axi_arvalid(ifu_arvalid), .s0_axi_arready(ifu_arready),
        .s0_axi_rdata(ifu_rdata),   .s0_axi_rvalid(ifu_rvalid),   .s0_axi_rready(ifu_rready),
        
        // Slave 1: LSU
        .s1_axi_awaddr(lsu_awaddr), .s1_axi_awvalid(lsu_awvalid), .s1_axi_awready(lsu_awready),
        .s1_axi_wdata(lsu_wdata_wire), .s1_axi_wstrb(lsu_wstrb), .s1_axi_wvalid(lsu_wvalid), .s1_axi_wready(lsu_wready),
        .s1_axi_bvalid(lsu_bvalid), .s1_axi_bready(lsu_bready),
        .s1_axi_araddr(lsu_araddr), .s1_axi_arvalid(lsu_arvalid), .s1_axi_arready(lsu_arready),
        .s1_axi_rdata(lsu_rdata_wire), .s1_axi_rvalid(lsu_rvalid), .s1_axi_rready(lsu_rready),
        
        // Master: Nối ra RAM
        .m_axi_awaddr(mem_awaddr), .m_axi_awvalid(mem_awvalid), .m_axi_awready(mem_awready),
        .m_axi_wdata(mem_wdata),   .m_axi_wstrb(mem_wstrb),     .m_axi_wvalid(mem_wvalid),   .m_axi_wready(mem_wready),
        .m_axi_bvalid(mem_bvalid), .m_axi_bready(mem_bready),
        .m_axi_araddr(mem_araddr), .m_axi_arvalid(mem_arvalid), .m_axi_arready(mem_arready),
        .m_axi_rdata(mem_rdata),   .m_axi_rvalid(mem_rvalid),   .m_axi_rready(mem_rready)
    );

    // 4. RAM (Mô hình bộ nhớ có độ trễ)
    axi4_ram_model #(
        .LATENCY(10),   // Giả lập độ trễ 10 chu kì
        .INIT_FILE("")  // Để trống, ta sẽ tự ghi dữ liệu
    ) DUT_RAM (
        .clk(clk), .rst_n(rst_n),
        .s_axi_awaddr(mem_awaddr), .s_axi_awvalid(mem_awvalid), .s_axi_awready(mem_awready),
        .s_axi_wdata(mem_wdata),   .s_axi_wstrb(mem_wstrb),     .s_axi_wvalid(mem_wvalid),   .s_axi_wready(mem_wready),
        .s_axi_bvalid(mem_bvalid), .s_axi_bready(mem_bready),
        .s_axi_araddr(mem_araddr), .s_axi_arvalid(mem_arvalid), .s_axi_arready(mem_arready),
        .s_axi_rdata(mem_rdata),   .s_axi_rvalid(mem_rvalid),   .s_axi_rready(mem_rready)
    );

    // =========================================================
    // TEST LOGIC
    // =========================================================
    
    // Clock Gen: 100MHz (Period 10ns)
    always #5 clk = ~clk;

    // Helper: Reset Pulse
    task apply_reset;
        begin
            rst_n = 0;
            #20;
            rst_n = 1;
            #20;
        end
    endtask

    // Helper: LSU Write
    task lsu_store_word(input [31:0] addr, input [31:0] data);
        begin
            @(posedge clk);
            lsu_we <= 1; lsu_re <= 0;
            lsu_mode <= 3'b010; // Word
            lsu_addr <= addr; lsu_wdata <= data;
            $display("[T=%0t] LSU REQ WRITE: Addr=%h, Data=%h", $time, addr, data);
            
            @(posedge clk);
            // Đợi hết stall (nghĩa là AXI done)
            while (lsu_stall) @(posedge clk);
            
            lsu_we <= 0; // Tắt lệnh
            $display("[T=%0t] LSU WRITE DONE", $time);
        end
    endtask

    // Helper: LSU Read
    task lsu_load_word(input [31:0] addr, input [31:0] expect_val);
        begin
            @(posedge clk);
            lsu_we <= 0; lsu_re <= 1;
            lsu_mode <= 3'b010; // Word
            lsu_addr <= addr;
            $display("[T=%0t] LSU REQ READ: Addr=%h", $time, addr);
            
            @(posedge clk);
            while (lsu_stall) @(posedge clk);
            
            lsu_re <= 0;
            #1; // Đợi ổn định để check
            if (lsu_rdata === expect_val)
                $display("[T=%0t] PASS: Read %h (Match)", $time, lsu_rdata);
            else
                $display("[T=%0t] FAIL: Read %h (Expected %h)", $time, lsu_rdata, expect_val);
        end
    endtask

    initial begin
        // Init signals
        clk = 0; rst_n = 0;
        pc = 32'h0;
        lsu_we=0; lsu_re=0; lsu_mode=0; lsu_addr=0; lsu_wdata=0;

        $display("=== START MEMORY SYSTEM TEST ===");
        apply_reset();

        // ----------------------------------------------------
        // TEST 1: Ghi dữ liệu vào RAM qua LSU
        // ----------------------------------------------------
        // Ghi số 0xDEADBEEF vào địa chỉ 0x100
        lsu_store_word(32'h00000100, 32'hDEADBEEF);
        
        #20;

        // ----------------------------------------------------
        // TEST 2: Đọc dữ liệu từ RAM qua LSU (Kiểm chứng Test 1)
        // ----------------------------------------------------
        lsu_load_word(32'h00000100, 32'hDEADBEEF);

        #20;

        // ----------------------------------------------------
        // TEST 3: Giả lập Fetch lệnh qua IFU
        // ----------------------------------------------------
        // Giả sử 0xDEADBEEF chính là mã lệnh ta vừa ghi
        $display("[T=%0t] IFU FETCH REQ: PC=0x100", $time);
        pc <= 32'h00000100; // Đổi PC
        
        @(posedge clk);
        // Đợi IFU Stall (đang đi lấy lệnh)
        while (ifu_stall) @(posedge clk);
        
        #1;
        if (instr === 32'hDEADBEEF)
            $display("[T=%0t] PASS: IFU Fetched %h (Match)", $time, instr);
        else
            $display("[T=%0t] FAIL: IFU Fetched %h (Expected DEADBEEF)", $time, instr);

        #20;

        // ----------------------------------------------------
        // TEST 4: Cache Hit Check
        // ----------------------------------------------------
        // Giữ nguyên PC, IFU sẽ không được Stall nữa (vì có cache)
        $display("[T=%0t] IFU CACHE CHECK (Same PC)", $time);
        @(posedge clk);
        if (ifu_stall == 0)
            $display("[PASS] IFU No Stall (Cache Hit works)");
        else
            $display("[FAIL] IFU Stalled again (Cache Missed?)");

        #20;

        // ----------------------------------------------------
        // TEST 5: Stress Test (Concurrent Access - Xung đột)
        // ----------------------------------------------------
        $display("[T=%0t] STRESS TEST: IFU Fetch & LSU Load same time", $time);
        // Thay đổi PC để IFU buộc phải miss -> Gọi AXI
        pc <= 32'h00000200; 
        
        // Đồng thời LSU gọi Load ở 0x100
        lsu_re <= 1; lsu_addr <= 32'h00000100;

        // Quan sát trên Waveform:
        // Interconnect sẽ cấp quyền cho LSU trước (vì ưu tiên cao hơn).
        // IFU sẽ bị Stall lâu hơn bình thường (đợi LSU xong mới đến lượt mình).
        
        repeat(50) @(posedge clk); // Chờ đủ lâu cho cả 2 xong
        lsu_re <= 0;

        $display("=== TEST FINISHED ===");
        $finish;
    end

endmodule